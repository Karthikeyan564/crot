`include "register_interface/typedef.svh"
`include "register_interface/assign.svh"

module mask_gen_top
    #(
      parameter int unsigned AXI_ADDR_WIDTH = 32,
      localparam int unsigned AXI_DATA_WIDTH = 32,
      parameter int unsigned AXI_ID_WIDTH,
      parameter int unsigned AXI_USER_WIDTH
      )
    (
     input logic clk_i,
     input logic rst_ni,
     input logic test_mode_i,

     AXI_BUS.Slave axi_slave
     );

    import mask_gen_reg_pkg::mask_gen_reg2hw_t;
    import mask_gen_reg_pkg::mask_gen_hw2reg_t;

    //Wiring Signals
    REG_BUS #(.ADDR_WIDTH(32), .DATA_WIDTH(32)) axi_to_regfile();
    mask_gen_reg2hw_t reg_file_to_ip;
    mask_gen_hw2reg_t ip_to_reg_file;

    axi_to_reg_intf #(
                      .ADDR_WIDTH(AXI_ADDR_WIDTH),
                      .DATA_WIDTH(AXI_DATA_WIDTH),
                      .ID_WIDTH(AXI_ID_WIDTH),
                      .USER_WIDTH(AXI_USER_WIDTH),
                      .DECOUPLE_W(0)
    ) i_axi2reg (
                 .clk_i,
                 .rst_ni,
                 .testmode_i(test_mode_i),
                 .in(axi_slave),
                 .reg_o(axi_to_regfile)
    );

    //Convert the REG_BUS interface to the struct signals used by autogenerated register file
    typedef logic [AXI_ADDR_WIDTH-1:0] addr_t;
    typedef logic [AXI_DATA_WIDTH-1:0] data_t;
    typedef logic [AXI_DATA_WIDTH/8-1:0] strb_t;
    `REG_BUS_TYPEDEF_REQ(reg_req_t, addr_t, data_t, strb_t);
    `REG_BUS_TYPEDEF_RSP(reg_rsp_t, data_t);
    reg_req_t to_reg_file_req;
    reg_rsp_t from_reg_file_rsp;

    `REG_BUS_ASSIGN_TO_REQ(to_reg_file_req, axi_to_regfile);
    `REG_BUS_ASSIGN_FROM_RSP(axi_to_regfile, from_reg_file_rsp);


    mask_gen_reg_top #(
    .reg_req_t(reg_req_t),
    .reg_rsp_t(reg_rsp_t)
    ) i_regfile (
                 .clk_i,
                 .rst_ni,
                 .devmode_i(1'b1),

                 //From the protocol converters to regfile
                 .reg_req_i(to_reg_file_req),
                 .reg_rsp_o(from_reg_file_rsp),

                 //Signals to mask gen IP
                 .reg2hw(reg_file_to_ip),
                 .hw2reg(ip_to_reg_file)
    );

    MGTop i_mask_gen (
                         .clk(clk_i),
                         .rst_n(rst_ni),
                         .clk_en(1'b1),
                         .pattern_w(reg_file_to_ip.mod_in.pattern_w.q),
			 .pattern(reg_file_to_ip.mod_in.pattern.q),
                         .repeatedPattern(reg_file_to_ip.mod_in.repeatedpattern.q),
                         .load_pattern(reg_file_to_ip.mod_in.load_pattern.q),
                         .mask_type(reg_file_to_ip.mod_in.mask_type.q),
                         .next(1'b1),//reg_file_to_ip.mod_in.next.q),
                         .imageResolution(reg_file_to_ip.mod_in.imgres.q),
                         .DOUT()//ip_to_reg_file.mod_out)
                         );

endmodule : mask_gen_top
